		
module adder_32bit(
  input  logic [31:0] A, B,
  input  logic        sel,      // 0: add, 1: sub (two's complement)
  output logic [31:0] OUT,
  output logic        CarryOut
);		
////////////////////////////////////////////////////////////////////////////		
//=============================
  // Tín hiệu nội bộ cho SPG
  //=============================
  logic [31:0] wb;        // B sau khi XOR với sel (đảo khi trừ)
  logic [31:0] G, P;      // Generate và Propagate từng bit
  logic [32:0] c;         // Carry tổng 33 bit (c[0] đến c[32])
		
    genvar i;

    generate
        for (i = 0; i < 32; i = i + 1) begin : SPG_block
            assign wb[i] = B[i] ^ sel;
            assign G[i] = A[i] & wb[i];
            assign P[i] = A[i] ^ wb[i];
            assign OUT[i] = P[i] ^ c[i];
        end
    endgenerate		
//=============================
// Gán liên kết carry tổng
//=============================
  	

 // Các nhóm P/G cho từng block 4-bit (Stage 1)
  //=============================
  logic P00, P01, P02, P03;  // nhóm 4-bit cho phần thấp
  logic G00, G01, G02, G03;
  logic P10, P11, P12, P13;  // nhóm 4-bit cho phần cao
  logic G10, G11, G12, G13;
 // Chia đôi 32-bit thành 2 nhóm 16-bit
  //=============================
  logic [15:0] c0, P0, G0;   // nhóm thấp (bit 0–15)
  logic [15:0] c1, P1, G1;   // nhóm cao  (bit 16–31)
  
  
// Carry-in cho từng nửa
  logic c0i, c1i;            // đầu vào của mỗi block
  assign c0i = sel;          // sel cũng chính là carry-in cho phép cộng/trừ	

//=============================
  // Liên kết dữ liệu 2 nửa
  //=============================
  assign P0 = P[15:0];
  assign G0 = G[15:0];
  assign P1 = P[31:16];
  assign G1 = G[31:16];

  //=============================	
  logic G20,P20,P21,G21;
  assign c = {c1, c0};
		
		
////////////////// c0LA_4bit staG0e 1 //////////// 
/////////////////					///////////
	assign c0[0] = c0i;
  assign c0[1] = G0[0] | (P0[0] & c0i);
  assign c0[2] = G0[1] | (P0[1] & G0[0]) | (P0[1] & P0[0] & c0i);
  assign c0[3] = G0[2] | (P0[2] & G0[1]) | (P0[2] & P0[1] & G0[0]) | (P0[2] & P0[1] & P0[0] & c0i);

  assign P00 =  P0[3]&P0[2]&P0[1]&P0[0];
  assign G00 = G0[3] | (P0[3] & G0[2]) | (P0[3] & P0[2] & G0[1]) | (P0[3] & P0[2] & P0[1] & G0[0]);
 

 ////////////////// c0LA_4bit staG0e 1 //////////// 
/////////////////					///////////
	
  assign c0[5] = G0[4] | (P0[4] & c0[4]);
  assign c0[6] = G0[5] | (P0[5] & G0[4]) | (P0[5] & P0[4] & c0[4]);
  assign c0[7] = G0[6] | (P0[6] & G0[5]) | (P0[6] & P0[5] & G0[4]) | (P0[6] & P0[5] & P0[4] & c0[4]);

  assign P01 = P0[7]&P0[6]&P0[5]&P0[4];
  assign G01 = G0[7] | (P0[7] & G0[6]) | (P0[7] & P0[6] & G0[5]) | (P0[7] & P0[6] & P0[5] & G0[4]);
 

 ////////////////// c0LA_4bit staG0e 1 //////////// 
/////////////////					///////////

  assign c0[9] = G0[8] | (P0[8] & c0[8]);
  assign c0[10] = G0[9] | (P0[9] & G0[8]) | (P0[9] & P0[8] & c0[8]);
  assign c0[11] = G0[10] | (P0[10] & G0[9]) | (P0[10] & P0[9] & G0[8]) | (P0[10] & P0[9] & P0[8] & c0[8]);

  assign P02 = P0[11]&P0[10]&P0[9]&P0[8];
  assign G02 = G0[11] | (P0[11] & G0[10]) | (P0[11] & P0[10] & G0[9]) | (P0[11] & P0[10] & P0[9] & G0[8]);
////////////////// c0LA_4bit staG0e 1 //////////// 
/////////////////					///////////

  assign c0[13] = G0[12] | (P0[12] & c0[12]);
  assign c0[14] = G0[13] | (P0[13] & G0[12]) | (P0[13] & P0[12] & c0[12]);
  assign c0[15] = G0[14] | (P0[14] & G0[13]) | (P0[14] & P0[13] & G0[12]) | (P0[14] & P0[13] & P0[12] & c0[12]);

  assign P03 = P0[15]&P0[14]&P0[13]&P0[12];
  assign G03 = G0[15] | (P0[15] & G0[14]) | (P0[15] & P0[14] & G0[13]) | (P0[15] & P0[14] & P0[13] & G0[12]);
  
  
  ////////////////// c0LA_4bit staG0e 2 //////////// 
/////////////////					///////////
  assign c0[4] = G00 | (P00 & c0i);
  assign c0[8] = G01 | (P01 & G00) | (P01 & P00 & c0i);
  assign c0[12] = G02 | (P02 & G01) | (P02 & P01 & G00) | (P02 & P01 & P00 & c0i);

  assign P20 =P03&P02&P01&P00;
  assign G20 = G03 | (P03 & G02) | (P03 & P02 & G01) | (P03 & P02 & P01 & G00);
  
  
  ////////////////////////// tang bit 16 dang sau//////////////////////////////////////////////////////////////////////
  ////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
  		
		
		
 
		
		
		
////////////////// c1LA_4bit staG1e 1 //////////// 
/////////////////					///////////
	assign c1[0] = c1i;
  assign c1[1] = G1[0] | (P1[0] & c1i);
  assign c1[2] = G1[1] | (P1[1] & G1[0]) | (P1[1] & P1[0] & c1i);
  assign c1[3] = G1[2] | (P1[2] & G1[1]) | (P1[2] & P1[1] & G1[0]) | (P1[2] & P1[1] & P1[0] & c1i);

  assign P10 =  P1[3]&P1[2]&P1[1]&P1[0];
  assign G10 = G1[3] | (P1[3] & G1[2]) | (P1[3] & P1[2] & G1[1]) | (P1[3] & P1[2] & P1[1] & G1[0]);
 

 ////////////////// c1LA_4bit staG1e 1 //////////// 
/////////////////					///////////
	
  assign c1[5] = G1[4] | (P1[4] & c1[4]);
  assign c1[6] = G1[5] | (P1[5] & G1[4]) | (P1[5] & P1[4] & c1[4]);
  assign c1[7] = G1[6] | (P1[6] & G1[5]) | (P1[6] & P1[5] & G1[4]) | (P1[6] & P1[5] & P1[4] & c1[4]);

  assign P11 = P1[7]&P1[6]&P1[5]&P1[4];
  assign G11 = G1[7] | (P1[7] & G1[6]) | (P1[7] & P1[6] & G1[5]) | (P1[7] & P1[6] & P1[5] & G1[4]);
 

 ////////////////// c1LA_4bit staG1e 1 //////////// 
/////////////////					///////////

  assign c1[9] = G1[8] | (P1[8] & c1[8]);
  assign c1[10] = G1[9] | (P1[9] & G1[8]) | (P1[9] & P1[8] & c1[8]);
  assign c1[11] = G1[10] | (P1[10] & G1[9]) | (P1[10] & P1[9] & G1[8]) | (P1[10] & P1[9] & P1[8] & c1[8]);

  assign P12 = P1[11]&P1[10]&P1[9]&P1[8];
  assign G12 = G1[11] | (P1[11] & G1[10]) | (P1[11] & P1[10] & G1[9]) | (P1[11] & P1[10] & P1[9] & G1[8]);
////////////////// c1LA_4bit staG1e 1 //////////// 
/////////////////					///////////

  assign c1[13] = G1[12] | (P1[12] & c1[12]);
  assign c1[14] = G1[13] | (P1[13] & G1[12]) | (P1[13] & P1[12] & c1[12]);
  assign c1[15] = G1[14] | (P1[14] & G1[13]) | (P1[14] & P1[13] & G1[12]) | (P1[14] & P1[13] & P1[12] & c1[12]);

  assign P13 = P1[15]&P1[14]&P1[13]&P1[12];
  assign G13 = G1[15] | (P1[15] & G1[14]) | (P1[15] & P1[14] & G1[13]) | (P1[15] & P1[14] & P1[13] & G1[12]);
  
  
  ////////////////// c1LA_4bit staG1e 2 //////////// 
/////////////////					///////////
  assign c1[4] = G10 | (P10 & c1i);
  assign c1[8] = G11 | (P11 & G10) | (P11 & P10 & c1i);
  assign c1[12] = G12 | (P12 & G11) | (P12 & P11 & G10) | (P12 & P11 & P10 & c1i);

  assign P21 =P13&P12&P11&P10 ;
  assign G21 = G13 | (P13 & G12) | (P13 & P12 & G11) | (P13 & P12 & P11 & G10);	
 




 
		
					///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
					/////////////////////////////////////////////// CLA 2bit ///////////////////////////////////////////////////////////////////////////////////////////////
					assign c1i = G20| (P20&c0i); 
					assign CarryOut = G21 | (P21 & G20)|(P21&P20&c0i);
					
					
	endmodule
	
					