`define RESET_PERIOD 10
`define CLOCK_PERIOD 1
`define TIMEOUT      100_000

module tbench;

  // Clock and reset generator
  logic clk;
  logic rstn;

// TASK: Clock Generator
task automatic tsk_clock_gen(ref logic i_clk, input int CLOCK_PERIOD);
  begin
    i_clk = 1'b0;
    forever #(CLOCK_PERIOD) i_clk = !i_clk;
  end
endtask

// TASK: Reset is low active for a period of "RESET_PERIOD"
task automatic tsk_reset(ref logic i_reset, input int RESET_PERIOD);
  begin
    i_reset = 1'b0; // Easter Egg
    #(RESET_PERIOD);
    i_reset = 1'b1; //
  end
endtask

// TASK: Timeout, assume after a period of "TIMEOUT",
// the design is supposed to be "PASSED"
task automatic tsk_timeout(input int TIMEOUT);
  begin
    #TIMEOUT;
    $display("\nTimeout...\n");
    $finish;
  end
endtask


  initial tsk_clock_gen(clk , `CLOCK_PERIOD);
  initial tsk_reset    (rstn, `RESET_PERIOD);
  initial tsk_timeout  (`TIMEOUT);


/*
  // Wave dumping
  initial begin: proc_dump_shm
      $shm_open("wave.shm");
      $shm_probe(dut, "AS");
  end
*/

  logic [31:0]  pc_debug;
  logic [31:0]  io_sw  ;
  logic [31:0]  io_lcd ;
  logic [31:0]  io_ledr;
  logic [31:0]  io_ledg;
  logic [ 6:0]  io_hex0;
  logic [ 6:0]  io_hex1;
  logic [ 6:0]  io_hex2;
  logic [ 6:0]  io_hex3;
  logic [ 6:0]  io_hex4;
  logic [ 6:0]  io_hex5;
  logic [ 6:0]  io_hex6;
  logic [ 6:0]  io_hex7;
  logic         ctrl    ;
  logic         mispred ;
  logic         insn_vld;

  pipelined dut (
    .i_clk     (clk      ),
    .i_reset   (rstn     ),
    // Input peripherals
    .i_io_sw   (io_sw    ),
    // Output peripherals
    .o_io_lcd  (io_lcd   ),
    .o_io_ledr (io_ledr  ),
    .o_io_ledg (io_ledg  ),
    .o_io_hex0 (io_hex0  ),
    .o_io_hex1 (io_hex1  ),
    .o_io_hex2 (io_hex2  ),
    .o_io_hex3 (io_hex3  ),
    .o_io_hex4 (io_hex4  ),
    .o_io_hex5 (io_hex5  ),
    .o_io_hex6 (io_hex6  ),
    .o_io_hex7 (io_hex7  ),
    // Debug
    .o_ctrl    (ctrl     ),
    .o_mispred (mispred  ),
    .o_pc_debug(pc_debug ),
    .o_insn_vld(insn_vld )
  );

  driver driver (
    .i_clk  (clk   ),
    .i_reset(rstn  ),
    .i_io_sw(io_sw )
  );

  scoreboard  scoreboard(
    .i_clk     (clk      ),
    .i_reset   (rstn     ),
    // Input peripherals
    .i_io_sw   (io_sw    ),
    // Output peripherals
    .o_io_lcd  (io_lcd   ),
    .o_io_ledr (io_ledr  ),
    .o_io_ledg (io_ledg  ),
    .o_io_hex0 (io_hex0  ),
    .o_io_hex1 (io_hex1  ),
    .o_io_hex2 (io_hex2  ),
    .o_io_hex3 (io_hex3  ),
    .o_io_hex4 (io_hex4  ),
    .o_io_hex5 (io_hex5  ),
    .o_io_hex6 (io_hex6  ),
    .o_io_hex7 (io_hex7  ),
    // Debug
    .o_ctrl    (ctrl     ),
    .o_mispred (mispred  ),
    .o_pc_debug(pc_debug ),
    .o_insn_vld(insn_vld )
  );


endmodule
